module rv32_decoder #()
  ();

endmodule
